`default_nettype none
`include "Router.svh"
`include "RouterPkg.pkg"

//////
////// Network on Chip (NoC) 18-341
////// Node module
//////
module Node #(parameter NODEID=0) (
    input  logic       clock, reset_n,

    input pkt_t        pkt_in,            // Data packet from TB
    input logic        pkt_in_avail,      // The packet from TB is available
    output logic       cQ_full,           // The queue is full

    output pkt_t       pkt_out,           // Outbound packet from node to TB
    output logic       pkt_out_avail,     // The oubound packet is available

    input logic        free_outbound,     // Node is free
    input logic        put_inbound,       // Node is transferring to router
    input logic [7:0]  payload_inbound,   // Data sent from node to router

    output logic       free_inbound,      // Router is free
    output logic       put_outbound,      // Router is transferring to node
    output logic [7:0] payload_outbound); // Data sent from node to router


endmodule : Node

/*
 *  Create a FIFO (First In First Out) buffer with depth 4 using the given
 *  interface and constraints
 *    - The buffer is initally empty
 *    - Reads are combinational, so data_out is valid unless empty is asserted
 *    - Removal from the queue is processed on the clock edge.
 *    - Writes are processed on the clock edge
 *    - If a write is pending while the buffer is full, do nothing
 *    - If a read is pending while the buffer is empty, do nothing
 */
module FIFO #(parameter WIDTH=32) (
    input logic              clock, reset_n,
    input logic [WIDTH-1:0]  data_in
    input logic              we, re
    output logic [WIDTH-1:0] data_out,
    output logic             full, empty);


endmodule : FIFO
